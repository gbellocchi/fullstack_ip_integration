module wide_alu_top
    `include "register_interface/typedef.svh"
    `include "register_interface/assign.svh"
    import wide_alu_reg_pkg::*;
    #(
        parameter int unsigned AXI_ADDR_WIDTH = 32,
        localparam int unsigned AXI_DATA_WIDTH = 32,
        parameter int unsigned AXI_ID_WIDTH = -1,
        parameter int unsigned AXI_USER_WIDTH = -1
    )(
        input logic                             clk_i,
        input logic                             rst_ni,
        input logic                             test_mode_i,
        AXI_BUS.Slave                           axi_in
    );

    REG_BUS axi_to_reg_file;

    axi_to_reg_intf #(
        parameter int ADDR_WIDTH = -1,
        parameter int DATA_WIDTH = -1,
        parameter int ID_WIDTH = -1,
        parameter int USER_WIDTH = -1,
        parameter bit DECOUPLE_W = 1
    ) axi_to_reg_intf_i (
        .clk_i,
        .rst_ni,
        .testmode_i,
        .in             ( axi_in            ),
        .reg_o          ( axi_to_reg_file   )
    );

    //Convert the REG_BUS interface to the struct signals used by the autogenerated interface
    typedef logic [AXI_DATA_WIDTH-1:0] data_t;
    typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
    typedef logic [AXI_DATA_WIDTH/8-1:0] strb_t;
    `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t)
    `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t)
    reg_req_t to_reg_file_req;
    reg_rsp_t from_reg_file_rsp;
    `REG_BUS_ASSIGN_TO_REQ(to_reg_file_req, axi_to_reg_file)
    `REG_BUS_ASSIGN_FROM_RSP(axi_to_reg_file, from_reg_file_rsp)

    wide_alu_reg2hw_t reg_file_to_ip;
    wide_alu_hw2reg_t ip_to_reg_file;

    wide_alu_reg_top  wide_alu_reg_top_i (
        .clk_i      ( clk_i             ),
        .rst_ni     ( rst_ni            ),
        .reg_req_i  ( to_reg_file_req   ),
        .reg_rsp_o  ( from_reg_file_rsp ),
        .reg2hw     ( reg_file_to_ip    ),
        .hw2reg     ( ip_to_reg_file    ), 
        .devmode_i  ( 1'b1              )
    );

    wide_alu i_wide_alu(
        .clk_i,
        .rst_ni,
        .trigger_i              ( reg_file_to_ip.ctrl1.trigger.q & reg_file_to_ip.ctrl1.trigger.qe      ),
        .clear_err_i            ( reg_file_to_ip.ctrl1.clear_err.q & reg_file_to_ip.ctrl1.clear_err.qe  ),
        .op_a_i                 ( reg_file_to_ip.op_a                                                   ),
        .op_b_i                 ( reg_file_to_ip.op_b                                                   ),
        .result_o               ( ip_to_reg_file.result                                                 ),
        .deaccel_factor_we_i    ( reg_file_to_ip.ctrl2.delay.qe                                         ),
        .deaccel_factor_i       ( reg_file_to_ip.ctrl2.delay.q                                          ),
        .deaccel_factor_o       ( ip_to_reg_file.ctrl2.delay.d                                          ),
        .op_sel_we_i            ( reg_file_to_ip.ctrl2.opsel.qe                                         ),
        .op_sel_i               ( wide_alu_pkg::optype_e'(reg_file_to_ip.ctrl2.opsel.q)                 ),
        .op_sel_o               ( wide_alu_pkg::optype_e'(ip_to_reg_file.ctrl2.opsel.d)                 ),
        .status_o               ( wide_alu_pkg::status_e'(ip_to_reg_file.status.d)                      )
    );